//  ###########################################################################
//
//  Licensed to the Apache Software Foundation (ASF) under one
//  or more contributor license agreements.  See the NOTICE file
//  distributed with this work for additional information
//  regarding copyright ownership.  The ASF licenses this file
//  to you under the Apache License, Version 2.0 (the
//  "License"); you may not use this file except in compliance
//  with the License.  You may obtain a copy of the License at
//
//  http://www.apache.org/licenses/LICENSE-2.0
//
//  Unless required by applicable law or agreed to in writing,
//  software distributed under the License is distributed on an
//  "AS IS" BASIS, WITHOUT WARRANTIES OR CONDITIONS OF ANY
//  KIND, either express or implied.  See the License for the
//  specific language governing permissions and limitations
//  under the License.
//
//  ###########################################################################

module top;
 
//------------------------------------------------------------------------------
//  Description:import package files
// -----------------------------------------------------------------------------   
  import uvm_pkg::*;
  
  initial
    begin
 //------------------------------------------------------------------------------
 //Description:setting the virtual interface and giving the name uart_iff
//------------------------------------------------------------------------------	    
	    uvm_config_db#(virtual uart_iff)::set(null,"*","VIF_0",if0);
//This will run the test class inside top	    
	    
	run_test();
    end
endmodule
  
